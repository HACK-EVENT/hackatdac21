/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 921;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00766564,
        64'h6e2c7663_73697200,
        64'h79746972_6f697270,
        64'h2d78616d_2c766373,
        64'h69720073_656d616e,
        64'h2d676572_00646564,
        64'h6e657478_652d7374,
        64'h70757272_65746e69,
        64'h00746669_68732d67,
        64'h65720073_74707572,
        64'h7265746e_6900746e,
        64'h65726170_2d747075,
        64'h72726574_6e690064,
        64'h65657073_2d746e65,
        64'h72727563_00736567,
        64'h6e617200_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h006c6564_6f6d0065,
        64'h6c626974_61706d6f,
        64'h6300736c_6c65632d,
        64'h657a6973_2300736c,
        64'h6c65632d_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'ha9000000_04000000,
        64'h03000000_01000000,
        64'h1d010000_04000000,
        64'h03000000_07000000,
        64'h0a010000_04000000,
        64'h03000000_00000004,
        64'h00000000_000010f1,
        64'hff000000_5b000000,
        64'h10000000_03000000,
        64'h09000000_02000000,
        64'h0b000000_02000000,
        64'hec000000_10000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00303030_30303131,
        64'h66666640_63696c70,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'h00010000_08000000,
        64'h03000000_00000c00,
        64'h00000000_000002f1,
        64'hff000000_5b000000,
        64'h10000000_03000000,
        64'h07000000_02000000,
        64'h03000000_02000000,
        64'hec000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000000_30303030,
        64'h32303166_66664074,
        64'h6e696c63_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_00010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h000000f1_ff000000,
        64'h5b000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_ec000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00303030,
        64'h30303031_66666640,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h00000000_e2000000,
        64'h04000000_03000000,
        64'h01000000_d7000000,
        64'h04000000_03000000,
        64'h01000000_c6000000,
        64'h04000000_03000000,
        64'h00c20100_b8000000,
        64'h04000000_03000000,
        64'ha0acb903_3f000000,
        64'h04000000_03000000,
        64'h00400d00_00000000,
        64'h00c0c2f0_ff000000,
        64'h5b000000_10000000,
        64'h03000000_00303535,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00303030_63326330,
        64'h66666640_74726175,
        64'h01000000_b1000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000000_01000000,
        64'h00000080_00000000,
        64'h5b000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_4f000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_a9000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_79000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_70000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_66000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h5f000000_05000000,
        64'h03000000_00000000,
        64'h5b000000_04000000,
        64'h03000000_00757063,
        64'h4f000000_04000000,
        64'h03000000_a0acb903,
        64'h3f000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h59730700_2c000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd4040000_28010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h0c050000_38000000,
        64'h34060000_edfe0dd0,
        64'h00000000_00000000,
        64'h000000ff_f0c2c004,
        64'h000000ff_f0c2c003,
        64'h000000ff_f0c2c001,
        64'h000000ff_f0c2c005,
        64'h28aed2a6_2b7e1516,
        64'h28aed2a6_2b7e1516,
        64'h09cf4f3c_abf71588,
        64'h28aed2a6_2b7e1516,
        64'h0ecd9fe8_d5761d02,
        64'h75836f93_a086fbf3,
        64'hc9d53cb7_c1a1ade9,
        64'he426e269_e2fcbb9f,
        64'h00000000_00000000,
        64'h2d2d2d2d_3c203032,
        64'h27636164_616b6361,
        64'h6820726f_6620646f,
        64'h6d206361_6d682074,
        64'h73657420_6f742065,
        64'h67617373_656d2065,
        64'h68742073_69207369,
        64'h6874203e_2d2d2d2d,
        64'h003afba2_1d24185b,
        64'hfc3fe2b0_10aefc11,
        64'h02a0edca_20ef2066,
        64'hb7d3585b_0f0fae19,
        64'h00000000_00000000,
        64'h00000000_00697261,
        64'h50206e69_206b6361,
        64'h6a207374_65656d20,
        64'h6d6f7472_6150206e,
        64'h69206b63_616a2073,
        64'h7465656d_206d6f74,
        64'h103cf58f_1d52a753,
        64'hc4029249_114f83c3,
        64'h35a2bdaa_77731ecd,
        64'habcf2236_cba76688,
        64'hc8ae6226_ab7d152f,
        64'hb03a0f32_413197af,
        64'ha8caf0fd_2245f678,
        64'h2266a7a6_5f44b551,
        64'h2ff23783_0024113a,
        64'h00000000_00000000,
        64'h0a0d216b_7020676e,
        64'h69726574_6e65202c,
        64'h656e6f64_20676e69,
        64'h64616f6c_206d6172,
        64'h00000000_0000000a,
        64'h00000a21_65726568,
        64'h20676e69_74736574,
        64'h000000ff_f5207000,
        64'h000000ff_f5203000,
        64'h000000ff_f5202000,
        64'h000000ff_f5209000,
        64'h000000ff_f5200000,
        64'h000000ff_f5208000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00008082_61457402,
        64'h70a2853e_4789c75f,
        64'hf0ef853e_fe944783,
        64'hc7fff0ef_853efe84,
        64'h4783dc7f_f0ef853e,
        64'h85bafdf4_4783fe84,
        64'h0713fcf4_0fa387aa,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853e47c1_fa07dbe3,
        64'h2781fec4_2783fef4,
        64'h262337fd_fec42783,
        64'hcc7ff0ef_853efe94,
        64'h4783cd1f_f0ef853e,
        64'hfe844783_e19ff0ef,
        64'h853e85ba_feb44783,
        64'hfe840713_fef405a3,
        64'h00f757b3_fd843703,
        64'h27810037_979bfec4,
        64'h2783a099_fef42623,
        64'h479dfca4_3c231800,
        64'hf022f406_71798082,
        64'h61457402_70a2853e,
        64'h47a1fa07_dae32781,
        64'hfec42783_fef42623,
        64'h37fdfec4_2783d35f,
        64'hf0ef853e_fe944783,
        64'hd3fff0ef_853efe84,
        64'h4783e87f_f0ef853e,
        64'h85bafeb4_4783fe84,
        64'h0713fef4_05a32781,
        64'h00f757bb_fdc42703,
        64'h27810037_979bfec4,
        64'h2783a0a1_fef42623,
        64'h478dfcf4_2e2387aa,
        64'h1800f022_f4067179,
        64'h80826121_744270e2,
        64'h853efec4_2783f607,
        64'hd3e32781_fe842783,
        64'hfef42423_37fdfe84,
        64'h2783fef4_26232785,
        64'hfec42783_db3ff0ef,
        64'h853efdf4_4783fcf4,
        64'h0fa30007_c78397ba,
        64'h16c78793_93011702,
        64'h00000797_0007871b,
        64'h8bbdfe04_2783fcf4,
        64'h2423fe84_278304f7,
        64'h70632781_fc842783,
        64'hfe842703_eb812781,
        64'hfe042783_fef42223,
        64'h02f757bb_47a9fe44,
        64'h2703fcf4_262340f7,
        64'h07bbfcc4_27032781,
        64'h02f707bb_fe442783,
        64'hfe042703_fef42023,
        64'h02f757bb_fe442783,
        64'hfcc42703_a859fef4,
        64'h242347a5_fef42223,
        64'ha007879b_3b9ad7b7,
        64'hfe042623_fcf42423,
        64'h87bafcf4_2623872e,
        64'h87aa0080_f822fc06,
        64'h71398082_61056462,
        64'h000100e7_8023fe04,
        64'h37830007_c70397ba,
        64'h21878793_00000797,
        64'h0007871b_8bbd2781,
        64'h0ff7f793_0047d79b,
        64'hfef44783_00e78023,
        64'h00074703_973623e7,
        64'h07130000_07170785,
        64'hfe043783_0007869b,
        64'h8bbd2781_fef44783,
        64'hfef407a3_feb43023,
        64'h87aa1000_ec221101,
        64'h80826145_740270a2,
        64'h853efec4_2783fbf9,
        64'h0007c783_fe043783,
        64'hfef42623_2785fec4,
        64'h2783fef4_30230785,
        64'hfe043783_ef3ff0ef,
        64'h853e0007_c783fe04,
        64'h3783a015_fef43023,
        64'hfd843783_fe042623,
        64'hfca43c23_1800f022,
        64'hf4067179_80826145,
        64'h740270a2_0001eb1f,
        64'hf0ef853e_02000593,
        64'h4907b783_00000797,
        64'hec3ff0ef_853e458d,
        64'h4987b783_00000797,
        64'hed3ff0ef_853e85ba,
        64'h4a07b783_00000797,
        64'h0ff7f713_27810087,
        64'hd79bfec4_2783ef1f,
        64'hf0ef00e7_951330b7,
        64'h879303ff_c7b785be,
        64'h0ff7f793_fec42783,
        64'hf0bff0ef_853e0800,
        64'h05934e27_b7830000,
        64'h0797f1df_f0ef853e,
        64'h45814ea7_b7830000,
        64'h0797fef4_262302f7,
        64'h57bbfdc4_27032781,
        64'h0047979b_fd842783,
        64'hfcf42c23_87bafcf4,
        64'h2e23872e_87aa1800,
        64'hf022f406_71798082,
        64'h61056442_60e20001,
        64'hf63ff0ef_00e79513,
        64'h30b78793_03ffc7b7,
        64'h85befef4_4783dfed,
        64'h87aafc7f_f0ef0001,
        64'hfef407a3_87aa1000,
        64'he822ec06_11018082,
        64'h01416402_60a2853e,
        64'h27810207_f7932781,
        64'h87aafd1f_f0ef853e,
        64'h5687b783_00000797,
        64'h0800e022_e4061141,
        64'h80826105_6462853e,
        64'h0ff7f793_0007c783,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61457422_000100e7,
        64'h8023fd74_4703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_0ba387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61217462,
        64'h853efd84_3783fce7,
        64'hece3fc84_3703fec4,
        64'h2783fef4_26232785,
        64'hfec42783_00e78023,
        64'h0ff77713_fd442703,
        64'h97bafd84_3703fec4,
        64'h2783a00d_fe042623,
        64'hfcf42a23_fcc43423,
        64'h87aefca4_3c230080,
        64'hfc227139_80826121,
        64'h7462853e_fd843783,
        64'hfce7e9e3_fc843703,
        64'hfec42783_fef42623,
        64'h2785fec4_2783c398,
        64'h431897b6_fd843683,
        64'h078afec4_2783973e,
        64'hfd043703_078afec4,
        64'h2783a025_fe042623,
        64'hfcc43423_fcb43823,
        64'hfca43c23_0080fc22,
        64'h71398082_61217462,
        64'h853efd84_3783fce7,
        64'he9e3fc84_3703fec4,
        64'h2783fef4_26232785,
        64'hfec42783_00e78023,
        64'h00074703_97b6fd84,
        64'h3683fec4_2783973e,
        64'hfd043703_fec42783,
        64'ha025fe04_2623fcc4,
        64'h3423fcb4_3823fca4,
        64'h3c230080_fc227139,
        64'h80826121_7462853e,
        64'hfec42783_fae7dfe3,
        64'h47850007_871bfe84,
        64'h2783fef4_24232785,
        64'hfe842783_fef42623,
        64'h4785a021_fe042623,
        64'h00f70563_8736439c,
        64'h97bafd04_3703078a,
        64'hfe842783_439497ba,
        64'hfd843703_078afe84,
        64'h2783a82d_fe042423,
        64'hfef42623_4785a8a1,
        64'h478100e7_f463fd04,
        64'h370397ba_fd043703,
        64'h078afcc4_2783a885,
        64'h478100e7_f463fd84,
        64'h370397ba_fd843703,
        64'h078afcc4_2783fcf4,
        64'h262387b2_fcb43823,
        64'hfca43c23_0080fc22,
        64'h71398082_61457422,
        64'h0001fef7_44e32781,
        64'h2701fdc4_2783fec4,
        64'h2703fef4_26232785,
        64'hfec42783_0001a039,
        64'hfe042623_fcf42e23,
        64'h87aa1800_f4227179,
        64'h80826161_640660a6,
        64'h0001f807_d8e32781,
        64'hfe442783_fef42223,
        64'h37fdfe44_2783fef4,
        64'h24232785_fe842783,
        64'he0bff0ef_fd843503,
        64'h85be863a_fec42703,
        64'h27812781_40f707bb,
        64'hfe842783_0007871b,
        64'h37fdfd44_2783eb8d,
        64'h27818b8d_fe442783,
        64'hfef42623_8fd98736,
        64'h27810007_c783fae4,
        64'h3c230017_8713fb84,
        64'h37830007_869b0087,
        64'h979bfec4_2783a0b5,
        64'hfef42223_37fdfc04,
        64'h2783fe04_2623fcf4,
        64'h2a234027_d79b9fb9,
        64'h01e7571b_41f7d71b,
        64'hfc042783_fe042423,
        64'hfcf43c23_97bafc84,
        64'h3703078e_fc446783,
        64'hfcf42023_87bafcf4,
        64'h22238736_fac43c23,
        64'h87aefca4_34230880,
        64'he0a2e486_715d8082,
        64'h61217442_70e20001,
        64'hfae7efe3_2781fec4,
        64'h2783fd04_2703fef4,
        64'h26232785_fec42783,
        64'hedbff0ef_fe043503,
        64'h85b6863e_439c97ba,
        64'hfc843703_078afec4,
        64'h67830007_869b37fd,
        64'h278140f7_07bbfec4,
        64'h2783fd04_2703a82d,
        64'hfe042623_fef43023,
        64'h97bafd84_3703078e,
        64'hfd446783_fcf42823,
        64'h87bafcf4_2a238736,
        64'hfcc43423_87aefca4,
        64'h3c230080_f822fc06,
        64'h71398082_616174e2,
        64'h640660a6_0001fae7,
        64'hece32781_fdc42783,
        64'hfc042703_fcf42e23,
        64'h2785fdc4_2783c09c,
        64'h278187aa_f37ff0ef,
        64'hfd043503_85befdc4,
        64'h278300f7_04b3fb84,
        64'h3703078a_93811782,
        64'h278137fd_278140f7,
        64'h07bbfdc4_2783fc04,
        64'h2703a081_fc042e23,
        64'hfcf43823_97bafc84,
        64'h3703078e_fc446783,
        64'hfcf42023_87bafcf4,
        64'h22238736_fac43c23,
        64'h87aefca4_34230880,
        64'hfc26e0a2_e486715d,
        64'h80826145_74220001,
        64'hc398fd04_2703fe84,
        64'h3783fef4_342397ba,
        64'hfd843703_078efd44,
        64'h6783fcf4_282387ba,
        64'hfcf42a23_873287ae,
        64'hfca43c23_1800f422,
        64'h71798082_61457422,
        64'h853e2781_439cfe84,
        64'h3783fef4_342397ba,
        64'hfd843703_078efd44,
        64'h6783fcf4_2a2387ae,
        64'hfca43c23_1800f422,
        64'h71798082_6129744a,
        64'h70ea853e_fe842783,
        64'hfef42423_87aa2a00,
        64'h00ef853e_85ba4621,
        64'hf6040793_f8040713,
        64'he29ff0ef_853e85ba,
        64'h8636fa04_0793f804,
        64'h0713fec4_26831380,
        64'h00ef853e_45e9863a,
        64'h46a1f404_07138be7,
        64'hb7830000_1797fe04,
        64'h2623f4f4_3c23f4e4,
        64'h3823f4d4_3423f4c4,
        64'h30236f9c_a4478793,
        64'h6b18a447_87136714,
        64'ha4478713_a447b603,
        64'h00001797_f6f43c23,
        64'hf6e43823_f6d43423,
        64'hf6c43023_6f9ca4e7,
        64'h87936b18_a4e78713,
        64'h6714a4e7_8713a4e7,
        64'hb6030000_1797fef4,
        64'h00230407_c783a687,
        64'h8793fce4_3c23fcd4,
        64'h3823fcc4_3423fcb4,
        64'h3023faa4_3c23fb04,
        64'h3823fb14_3423fa64,
        64'h30237f18_a6878713,
        64'h7b14a687_87137710,
        64'ha6878713_730ca687,
        64'h87136f08_a6878713,
        64'h01073803_a6878713,
        64'h00873883_a6878713,
        64'ha687b303_00001797,
        64'h0180f922_fd067131,
        64'h80826121_744270e2,
        64'h853e4781_190000ef,
        64'h853e45c9_fd043603,
        64'h46a19a27_b7830000,
        64'h1797d3fd_278187aa,
        64'h142000ef_853e45c5,
        64'h9b87b783_00001797,
        64'h3a4000ef_4511a021,
        64'h3ac000ef_45511900,
        64'h00ef853e_45814601,
        64'h9d87b783_00001797,
        64'h1a2000ef_853e4581,
        64'h46059ea7_b7830000,
        64'h1797a01d_1b6000ef,
        64'h853e4581_46119fe7,
        64'hb7830000_17971c80,
        64'h00ef853e_45814615,
        64'ha107b783_00001797,
        64'hc7852781_fcc42783,
        64'h32e000ef_853e4585,
        64'hfd843603_04000693,
        64'ha307b783_00001797,
        64'hd3fd2781_87aa1d00,
        64'h00ef853e_4581a467,
        64'hb7830000_17974320,
        64'h00ef4505_a021fef4,
        64'h3423fd84_3783fcf4,
        64'h262387b2_fcb43823,
        64'hfca43c23_0080f822,
        64'hfc067139_80826149,
        64'h640a60aa_853efec4,
        64'h2783fef4_262387aa,
        64'h4a2000ef_853e85ba,
        64'h4621f784_0793f984,
        64'h0713bd3f_f0ef853e,
        64'h85bafb84_0793f984,
        64'h0713f8f4_3823f8e4,
        64'h3423f8d4_3023f6c4,
        64'h3c236f9c_b9c78793,
        64'h6b18b9c7_87136714,
        64'hb9c78713_b9c7b603,
        64'h00001797_fe041423,
        64'hfe042223_fef42023,
        64'h579cbaa7_8793fce4,
        64'h3c23fcd4_3823fcc4,
        64'h3423fcb4_3023faa4,
        64'h3c237318_baa78713,
        64'h6f14baa7_87136b10,
        64'hbaa78713_670cbaa7,
        64'h8713baa7_b5030000,
        64'h17970900_e122e506,
        64'h71758082_61217462,
        64'h853e2781_4037d79b,
        64'h9fb901d7_571b41f7,
        64'hd71bfe44_2783f6e7,
        64'hc0e32781_fec42783,
        64'h0007871b_27a1fdc4,
        64'h2783fef4_26232785,
        64'hfec42783_00078023,
        64'h97bafc04_3703fec4,
        64'h2783a801_00e78023,
        64'h0ff6f713_97bafc04,
        64'h3703fec4_278300f7,
        64'h56b3fc84_3703fd44,
        64'h6783fcf4_2a230037,
        64'h979b2781_40f707bb,
        64'hfd842783_471dfcf4,
        64'h2c2340f7_07bbfdc4,
        64'h2783fec4_270304f7,
        64'h44632781_2701fdc4,
        64'h2783fec4_2703a095,
        64'h00e78023_f8000713,
        64'h97bafc04_3703fec4,
        64'h278300f7_1c632781,
        64'h2701fe04_2783fec4,
        64'h2703a849_fef42623,
        64'hfe042783_fcf42e23,
        64'h9fb9fe04_27032781,
        64'h37e12781_4037d79b,
        64'h9fb901d7_571b41f7,
        64'hd71bfe44_2783fef4,
        64'h20234037_d79b9fb9,
        64'h01d7571b_41f7d71b,
        64'hfe842783_fef42223,
        64'h278140f7_07bbfe84,
        64'h27832000_0713a801,
        64'h278140f7_07bbfe84,
        64'h27834000_071300e7,
        64'hda631c00_07930007,
        64'h871bfe84_2783fef4,
        64'h24231ff7_f7932781,
        64'hfc843783_fcb43023,
        64'hfca43423_0080fc22,
        64'h71398082_44010113,
        64'h43013403_43813083,
        64'h853e4781_480000ef,
        64'h853e45c9_bc043603,
        64'h46a1c8a7_b7830000,
        64'h1797de07_8de32781,
        64'hfec42783_d3fd2781,
        64'h87aa43c0_00ef853e,
        64'h45c5caa7_b7830000,
        64'h179769e0_00ef4511,
        64'ha0216a60_00ef4551,
        64'h48a000ef_853e4581,
        64'h4601cca7_b7830000,
        64'h179749c0_00ef853e,
        64'h45814609_cdc7b783,
        64'h00001797_576000ef,
        64'h853a4585_863e46c1,
        64'h04078793_bd040793,
        64'hcf87b703_00001797,
        64'hd3fd2781_87aa4a00,
        64'h00ef853e_4581d0e7,
        64'hb7830000_17977020,
        64'h00ef4505_a02108e7,
        64'hd3630400_07930007,
        64'h871bfd04_2783d3fd,
        64'h278187aa_4ce000ef,
        64'h853e45c5_d3c7b783,
        64'h00001797_730000ef,
        64'h4511a021_738000ef,
        64'h455151c0_00ef853e,
        64'h45814601_d5c7b783,
        64'h00001797_52e000ef,
        64'h853e4581_4609d6e7,
        64'hb7830000_1797a01d,
        64'hfe042423_546000ef,
        64'h853e4581_4601d867,
        64'hb7830000_17975580,
        64'h00ef853e_45814605,
        64'hd987b783_00001797,
        64'hc7952781_fe842783,
        64'h6be000ef_853e4585,
        64'h863a0400_0693bd04,
        64'h0713dba7_b7830000,
        64'h1797d3fd_278187aa,
        64'h562000ef_853e4581,
        64'hdd07b783_00001797,
        64'h7c4000ef_4505a021,
        64'hfcf42823_87aa1800,
        64'h00ef853a_85bebd04,
        64'h0793873e_27810037,
        64'h979bfe44_2783c785,
        64'h2781fec4_2783fc04,
        64'h2823fae7_d7e303f0,
        64'h07930007_871bfd44,
        64'h2783fef4_22232785,
        64'hfe442783_fcf42a23,
        64'h2785fd44_278300e7,
        64'h80230007_4703fcd4,
        64'h3c230017_8693fd84,
        64'h3783bcf4_34230017,
        64'h0793bc84_3703a099,
        64'hfef42623_4785e789,
        64'h0007c783_bc843783,
        64'ha0a1fc04_2a23fcf4,
        64'h3c23bd04_0793fce7,
        64'hdee307f0_07930007,
        64'h871bfe04_2783fef4,
        64'h20232785_fe042783,
        64'hbe078023_97baff04,
        64'h0713fe04_2783a829,
        64'hfe042023_a409fe04,
        64'h2223fef4_24234785,
        64'hfe042623_bcb43023,
        64'hbca43423_44010413,
        64'h42813823_42113c23,
        64'hbc010113_80826165,
        64'h740670a6_853efe84,
        64'h2783fef4_242387aa,
        64'h0fb000ef_853e85ba,
        64'h4611f904_0793fa04,
        64'h0713e75f_f0ef853e,
        64'h85bafd84_0793fc84,
        64'h0713fa04_0613fec4,
        64'h26837940_00ef853e,
        64'h4595863a_4699fb04,
        64'h0713f027_b7830000,
        64'h1797fe04_2623f8f4,
        64'h3c23679c_fbc78793,
        64'hf8e43823_fbc7b703,
        64'h00001797_fcf43023,
        64'h6b9cfc47_8793fae4,
        64'h3c236718_fc478713,
        64'hfae43823_fc47b703,
        64'h00001797_fcf43823,
        64'h679cfca7_8793fce4,
        64'h3423fca7_b7030000,
        64'h1797fef4_3023679c,
        64'hfd078793_fce43c23,
        64'hfd07b703_00001797,
        64'h1880f0a2_f4867159,
        64'h80826145_740270a2,
        64'h853e4781_798000ef,
        64'h853e45b1_fd843603,
        64'h4691f927_b7830000,
        64'h1797d3fd_278187aa,
        64'h74a000ef_853e45ad,
        64'hfa87b783_00001797,
        64'h1ad000ef_4511a021,
        64'h792000ef_853e4581,
        64'h4601fc27_b7830000,
        64'h1797d3fd_278187aa,
        64'h77a000ef_853e4581,
        64'hfd87b783_00001797,
        64'h1dd000ef_4505a021,
        64'h7c2000ef_853e4581,
        64'h4605ff27_b7830000,
        64'h17977d40_00ef853e,
        64'h45814601_0047b783,
        64'h00001797_0af000ef,
        64'h853e45c1_fe043603,
        64'h469101a7_b7830000,
        64'h17970c50_00ef853e,
        64'h4585fe84_36034691,
        64'h0307b783_00001797,
        64'h013000ef_853e0200,
        64'h0593863a_fd442703,
        64'h0487b783_00001797,
        64'hfcf42a23_87b6fcc4,
        64'h3c23feb4_3023fea4,
        64'h34231800_f022f406,
        64'h71798082_01416402,
        64'h60a2853e_4781a011,
        64'h478500f7_14634785,
        64'h873e87aa_fa1ff0ef,
        64'h0800e022_e4061141,
        64'h80826105_644260e2,
        64'h853e4785_d3f12781,
        64'h87aa04d0_00ef853e,
        64'h45b90a27_b7830000,
        64'h1797a829_478100e7,
        64'hd4636807_87930098,
        64'h97b70007_871bfec4,
        64'h2783fef4_26232785,
        64'hfec42783_2d1000ef,
        64'h4505a02d_fe042623,
        64'h1000e822_ec061101,
        64'h80822601_01132481,
        64'h34832501_34032581,
        64'h3083853e_4781a011,
        64'h47810050_0293c63f,
        64'hf0efe399_2781fc04,
        64'h2783c789_2781fc44,
        64'h2783cb89_2781fc84,
        64'h2783cf89_2781fd04,
        64'h2783c38d_2781fd44,
        64'h2783fcf4_2023fbc4,
        64'h2783faf4_2e2387aa,
        64'h0b4000ef_fcf42223,
        64'hfbc42783_fcf42423,
        64'hfbc42783_fcf42a23,
        64'hfbc42783_faf42e23,
        64'h4785fcf4_20234785,
        64'hfcf42223_4785fcf4,
        64'h24234785_fcf42623,
        64'h4785fcf4_28234785,
        64'hfcf42a23_47856b70,
        64'h00ef1ca5_05130000,
        64'h15176c30_00ef1ce5,
        64'h05130000_15170d40,
        64'h10ef853e_639cfce4,
        64'h3c230087_8713fd84,
        64'h37830e80_10ef853e,
        64'hfd843783_6ed000ef,
        64'h1f850513_00001517,
        64'h0fe010ef_853e639c,
        64'hfce43c23_00878713,
        64'hfd843783_112010ef,
        64'h853efd84_3783fcf4,
        64'h3c230792_12978793,
        64'h080017b7_725000ef,
        64'h23050513_00001517,
        64'h136010ef_853e639c,
        64'hfce43c23_00878713,
        64'hfd843783_14a010ef,
        64'h853efd84_378374f0,
        64'h00ef25a5_05130000,
        64'h15171600_10ef853e,
        64'h639cfce4_3c230087,
        64'h8713fd84_37831740,
        64'h10ef853e_fd843783,
        64'hfcf43c23_07fe4785,
        64'h781000ef_27c50513,
        64'h00001517_6db000ef,
        64'hca078513_03b9b7b7,
        64'h20078593_67f11607,
        64'h9a632781_87aadebf,
        64'hf0efb525_257000ef,
        64'h853e459d_46012a67,
        64'hb7830000_17972690,
        64'h00ef853e_45994605,
        64'h2b87b783_00001797,
        64'h5cb000ef_853e85ba,
        64'h8636da04_0713fa44,
        64'h6683fa84_3783cf81,
        64'h2781fb84_27835e90,
        64'h00ef853e_85ba8636,
        64'hda040793_fa446683,
        64'hfb043703_cf812781,
        64'hfb842783_faf42223,
        64'h87aa28d0_00ef853e,
        64'h458530a7_b7830000,
        64'h1797faf4_34238fc5,
        64'h93811782_278187aa,
        64'h2ab000ef_853e4591,
        64'h3287b783_00001797,
        64'h02079493_fa843783,
        64'hfaf43423_93811782,
        64'h278187aa_2cf000ef,
        64'h853e4595_34c7b783,
        64'h00001797_faf43823,
        64'h8fc59381_17822781,
        64'h87aa2ed0_00ef853e,
        64'h458936a7_b7830000,
        64'h17970207_9493fb04,
        64'h3783faf4_38239381,
        64'h17822781_87aa3110,
        64'h00ef853e_458d38e7,
        64'hb7830000_17970001,
        64'hbff15770_00ef4515,
        64'he7892781_fb842783,
        64'hfaf42c23_87aa3390,
        64'h00ef853e_45a53b67,
        64'hb7830000_17973790,
        64'h00ef853e_45814601,
        64'h3c87b783_00001797,
        64'hfcf718e3_4791873e,
        64'h278187aa_367000ef,
        64'h853e459d_3e47b783,
        64'h00001797_3a7000ef,
        64'h853e459d_46113f67,
        64'hb7830000_17975db0,
        64'h00ef4515_a8293c10,
        64'h00ef853e_459d4611,
        64'h4107b783_00001797,
        64'hd3f92781_87aa3a90,
        64'h00ef853e_45814267,
        64'hb7830000_179760b0,
        64'h00ef453d_f71ff0ef,
        64'h00f71463_4785873e,
        64'h278187aa_3cf000ef,
        64'h853e45a1_44c7b783,
        64'h00001797_ae2d4781,
        64'h02f71763_4785873e,
        64'h278187aa_3ef000ef,
        64'h853e45a1_46c7b783,
        64'h00001797_1cf71f63,
        64'h4785873e_278187aa,
        64'hfd5ff0ef_14802491,
        64'h34232481_38232411,
        64'h3c23da01_01138082,
        64'h61056462_853efec4,
        64'h2783fef4_2623f140,
        64'h27f31000_ec221101,
        64'h00000000_ffdff06f,
        64'h10500073_65458593,
        64'h00001597_f1402573,
        64'h00048067_01f49493,
        64'h0010049b_66c58593,
        64'h00001597_f1402573,
        64'h04e000ef_00410133,
        64'h00a11133_01111113,
        64'h00100113_f1402573,
        64'h01f21213_00100213
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
