/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom_linux (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 682;

    const logic [RomSize-1:0][63:0] mem = {
        64'h000000ff_f0c2c004,
        64'h000000ff_f0c2c003,
        64'h000000ff_f0c2c001,
        64'h000000ff_f0c2c005,
        64'h00000000_000a0d31,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_00000000,
        64'h2d2d2d2d_3c203032,
        64'h27636164_616b6361,
        64'h6820726f_6620646f,
        64'h6d206361_6d682074,
        64'h73657420_6f742065,
        64'h67617373_656d2065,
        64'h68742073_69207369,
        64'h6874203e_2d2d2d2d,
        64'h00000000_00766564,
        64'h6e2c7663_73697200,
        64'h79746972_6f697270,
        64'h2d78616d_2c766373,
        64'h69720073_656d616e,
        64'h2d676572_00646564,
        64'h6e657478_652d7374,
        64'h70757272_65746e69,
        64'h00746669_68732d67,
        64'h65720073_74707572,
        64'h7265746e_6900746e,
        64'h65726170_2d747075,
        64'h72726574_6e690064,
        64'h65657073_2d746e65,
        64'h72727563_00736567,
        64'h6e617200_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h006c6564_6f6d0065,
        64'h6c626974_61706d6f,
        64'h6300736c_6c65632d,
        64'h657a6973_2300736c,
        64'h6c65632d_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'ha9000000_04000000,
        64'h03000000_01000000,
        64'h1d010000_04000000,
        64'h03000000_07000000,
        64'h0a010000_04000000,
        64'h03000000_00000004,
        64'h00000000_000010f1,
        64'hff000000_5b000000,
        64'h10000000_03000000,
        64'h09000000_02000000,
        64'h0b000000_02000000,
        64'hec000000_10000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00303030_30303131,
        64'h66666640_63696c70,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'h00010000_08000000,
        64'h03000000_00000c00,
        64'h00000000_000002f1,
        64'hff000000_5b000000,
        64'h10000000_03000000,
        64'h07000000_02000000,
        64'h03000000_02000000,
        64'hec000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000000_30303030,
        64'h32303166_66664074,
        64'h6e696c63_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_00010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h000000f1_ff000000,
        64'h5b000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_ec000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00303030,
        64'h30303031_66666640,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h00000000_e2000000,
        64'h04000000_03000000,
        64'h01000000_d7000000,
        64'h04000000_03000000,
        64'h01000000_c6000000,
        64'h04000000_03000000,
        64'h00c20100_b8000000,
        64'h04000000_03000000,
        64'ha0acb903_3f000000,
        64'h04000000_03000000,
        64'h00400d00_00000000,
        64'h00c0c2f0_ff000000,
        64'h5b000000_10000000,
        64'h03000000_00303535,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00303030_63326330,
        64'h66666640_74726175,
        64'h01000000_b1000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000000_01000000,
        64'h00000080_00000000,
        64'h5b000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_4f000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_a9000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_79000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_70000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_66000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h5f000000_05000000,
        64'h03000000_00000000,
        64'h5b000000_04000000,
        64'h03000000_00757063,
        64'h4f000000_04000000,
        64'h03000000_a0acb903,
        64'h3f000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h59730700_2c000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd4040000_28010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h0c050000_38000000,
        64'h34060000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000a0d,
        64'h0a0d0a0d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_0a0d2020,
        64'h20202020_20202020,
        64'h34202f20_426b2034,
        64'h36202020_3a636f73,
        64'h7341202f_20657a69,
        64'h53202032_4c0a0d20,
        64'h20202020_20202020,
        64'h2034202f_20426b20,
        64'h38202020_203a636f,
        64'h73734120_2f20657a,
        64'h69532035_314c0a0d,
        64'h20202020_20202020,
        64'h20203420_2f20426b,
        64'h20382020_20203a63,
        64'h6f737341_202f2065,
        64'h7a695320_44314c0a,
        64'h0d202020_20202020,
        64'h20202034_202f2042,
        64'h6b203631_2020203a,
        64'h636f7373_41202f20,
        64'h657a6953_2049314c,
        64'h0a0d2020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20200a0d_20202020,
        64'h20202020_20202020,
        64'h20202020_424d2036,
        64'h39303420_20202020,
        64'h20202020_3a657a69,
        64'h53204d41_52440a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202067_69666e6f,
        64'h635f6873_656d6432,
        64'h20202020_20202020,
        64'h2020203a_6b726f77,
        64'h74654e0a_0d202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h7a484d20_32362020,
        64'h20202020_2020203a,
        64'h71657246_2065726f,
        64'h430a0d20_20202020,
        64'h20202020_20202020,
        64'h20202020_20203120,
        64'h20202020_20202020,
        64'h2020203a_7365726f,
        64'h43230a0d_20202020,
        64'h20202020_20202020,
        64'h20202020_20202031,
        64'h20202020_20202020,
        64'h20203a73_656c6954,
        64'h2d59230a_0d202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h31202020_20202020,
        64'h2020203a_73656c69,
        64'h542d5823_0a0d2020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20200a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202035_313a3330,
        64'h3a303220_31323032,
        64'h20303120_67754120,
        64'h20202020_2020203a,
        64'h65746144_20646c69,
        64'h75420a0d_20202020,
        64'h20202020_20202020,
        64'h20202020_20202031,
        64'h66202020_20202020,
        64'h203a6472_616f4220,
        64'h41475046_0a0d2020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20200a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202032_62313565,
        64'h33653020_2020203a,
        64'h6e6f6973_72655620,
        64'h656e6169_72410a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202032_62313565,
        64'h33653020_3a6e6f69,
        64'h73726556_206e6f74,
        64'h69506e65_704f0a0d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h0a0d2d2d_20202020,
        64'h20206d72_6f667461,
        64'h6c502065_6e616972,
        64'h412b6e6f_7469506e,
        64'h65704f20_20202020,
        64'h2d2d0a0d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_0a0d0a0d,
        64'h28aed2a6_2b7e1516,
        64'h28aed2a6_2b7e1516,
        64'h09cf4f3c_abf71588,
        64'h28aed2a6_2b7e1516,
        64'h0ecd9fe8_d5761d02,
        64'h75836f93_a086fbf3,
        64'hc9d53cb7_c1a1ade9,
        64'he426e269_e2fcbb9f,
        64'h003afba2_1d24185b,
        64'hfc3fe2b0_10aefc11,
        64'h02a0edca_20ef2066,
        64'hb7d3585b_0f0fae19,
        64'h00000000_00000000,
        64'h00000000_00697261,
        64'h50206e69_206b6361,
        64'h6a207374_65656d20,
        64'h6d6f7472_6150206e,
        64'h69206b63_616a2073,
        64'h7465656d_206d6f74,
        64'h103cf58f_1d52a753,
        64'hc4029249_114f83c3,
        64'h35a2bdaa_77731ecd,
        64'habcf2236_cba76688,
        64'hc8ae6226_ab7d152f,
        64'hb03a0f32_413197af,
        64'ha8caf0fd_2245f678,
        64'h2266a7a6_5f44b551,
        64'h2ff23783_0024113a,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h000000ff_f5208000,
        64'h000000ff_f5200000,
        64'h000000ff_f5209000,
        64'h000000ff_f5202000,
        64'h000000ff_f5203000,
        64'h000000ff_f5207000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_80826105,
        64'h450164a2_644260e2,
        64'h00500293_fa5ff0ef,
        64'he119c011_c0999b1f,
        64'hf0ef842a_cf9ff0ef,
        64'h84aaa5df_f0efe55f,
        64'hf0efc9a5_05130000,
        64'h1517e61f_f0efc8e5,
        64'h05130000_1517e13f,
        64'hf0efe426_e822ec06,
        64'hca050513_20058593,
        64'h110103b9_b53765f1,
        64'hffdff06f_10500073,
        64'h63858593_00000597,
        64'hf1402573_80826105,
        64'h450960e2_e27ff0ef,
        64'h00914503_e2fff0ef,
        64'h00814503_eddff0ef,
        64'hec06002c_11018082,
        64'h61454541_694264e2,
        64'h740270a2_fe9410e3,
        64'he53ff0ef_00914503,
        64'he5bff0ef_34610081,
        64'h4503f0bf_f0ef0ff5,
        64'h7513002c_00895533,
        64'h54e10380_0413892a,
        64'hf406e84a_ec26f022,
        64'h71798082_61454521,
        64'h694264e2_740270a2,
        64'hfe9410e3_e97ff0ef,
        64'h00914503_e9fff0ef,
        64'h34610081_4503f4ff,
        64'hf0ef0ff5_7513002c,
        64'h0089553b_54e14461,
        64'h892af406_e84aec26,
        64'hf0227179_80826121,
        64'h6b026aa2_6a4269e2,
        64'h790274a2_854e7442,
        64'h70e2fd59_14e30004,
        64'h851b397d_85d2ee9f,
        64'hf0ef2985_0007c503,
        64'h97ba18c7_87938b3d,
        64'h00000797_00ba7e63,
        64'he3990364_543b0285,
        64'h74bb0007_079b0009,
        64'h0a1b0285_573b5afd,
        64'h4b294981_4925a004,
        64'h0413e852_f426fc06,
        64'he05ae456_ec4ef04a,
        64'h3b9ad437_f8227139,
        64'h808200f5_80230007,
        64'hc78300e5_80a397aa,
        64'h81110007_4703973e,
        64'h00f57713_1ec78793,
        64'h00000797_b7d50405,
        64'hf63ff0ef_853e8082,
        64'h610564a2_644260e2,
        64'he7914094_053b0004,
        64'h4783842a_84aaec06,
        64'he426e822_11018082,
        64'h00e78023_02000713,
        64'he707b783_00001797,
        64'h00f70023_478d00a6,
        64'h80230ff5_751300c7,
        64'h80230085_551b0ff5,
        64'h761307ba_30b78793,
        64'h03ffc7b7_00f70023,
        64'hf8000793_00068023,
        64'hea07b703_00001797,
        64'hea07b683_00001797,
        64'h02b5553b_0045959b,
        64'h808200a7_802307ba,
        64'h30b78793_03ffc7b7,
        64'hdbe50207_f7930007,
        64'hc783ec27_b7830000,
        64'h17978082_02057513,
        64'h0007c503_ed47b783,
        64'h00001797_80820005,
        64'h45038082_00b50023,
        64'h8082bfd5_078500b7,
        64'h80238082_00c79363,
        64'h962a87aa_bfc5fee7,
        64'hae230591_07914198,
        64'h808200c5_9363962e,
        64'h87aa060a_b7fdfee7,
        64'h8fa30585_07850005,
        64'hc7038082_00c59363,
        64'h962e87aa_80824501,
        64'hafdff06f_00064463,
        64'h80826129_744a70ea,
        64'hb0dff0ef_1028002c,
        64'hf25ff0ef_10a84601,
        64'h002cbcdf_f0ef45e9,
        64'h00b046a1_3447b503,
        64'h00000797_03c000ef,
        64'h00a80200_06130c04,
        64'h059304a0_00ef1028,
        64'h02000613_0a040593,
        64'h058000ef_45640413,
        64'hfd060000_041710a8,
        64'hf2e58593_04100613,
        64'hf9220000_15977131,
        64'hbf654511_bf6d0007,
        64'ha023c398_47053967,
        64'hb7830000_0797b745,
        64'hc9bff0ef_45058082,
        64'h61054501_690264a2,
        64'h644260e2_c25ff0ef,
        64'h45c946a1_8622cb95,
        64'h27810885_27833c67,
        64'hb5030000_0797cc9f,
        64'hf0ef4551_c3984711,
        64'hc3984715_3dc7b783,
        64'h00000797_c4a1c9ff,
        64'hf0ef4585_864a0400,
        64'h0693c7b9_2781411c,
        64'h3f87b503_00000797,
        64'h84b2842e_892aec06,
        64'he04ae426_e8221101,
        64'h80826149_640a60aa,
        64'hbfdff0ef_1028002c,
        64'he5bff0ef_00a8002c,
        64'h118000ef_06011c23,
        64'hda821028_08040593,
        64'h02000613_12c000ef,
        64'he50600a8_02c00613,
        64'h04840593_53440413,
        64'h00000417_e1227175,
        64'hbdf54b85_8c2ac4ff,
        64'hf0ef858a_0034951b,
        64'hb7ed4511_ffb12781,
        64'h0887a783_47c7b783,
        64'h00000797_d77ff0ef,
        64'h0007a023_0137a023,
        64'h45514927_b7830000,
        64'h0797d25f_f0ef4585,
        64'h009046c1_d7fd2781,
        64'h411c4aa7_b5030000,
        64'h0797da5f_f0ef4505,
        64'hb7514511_b7490137,
        64'ha0234c27_b7830000,
        64'h0797b79d_dbfff0ef,
        64'h45058082_45010113,
        64'h45014001_3c034081,
        64'h3b834101_3b034181,
        64'h3a834201_3a034281,
        64'h39834301_39034381,
        64'h34834401_34034481,
        64'h3083d6bf_f0ef45c9,
        64'h46a18652_50c7b503,
        64'h00000797_f80b81e3,
        64'h895e0787_c6630400,
        64'h0793c7a5_27810887,
        64'ha78352a7_b7830000,
        64'h0797e25f_f0ef4551,
        64'h0007a023_0167a023,
        64'h5407b783_00000797,
        64'h08090163_dfdff0ef,
        64'h4585860a_04000693,
        64'hc7c12781_411c55e7,
        64'hb5030000_07974c01,
        64'h4b81fe86_97e30785,
        64'h24850405_00e78023,
        64'h10070663_00044703,
        64'h04040693_878aff57,
        64'h9be30785_00070023,
        64'h00f10733_47814b05,
        64'h49890800_0a934905,
        64'h44818a2e_842a4181,
        64'h30234171_34234411,
        64'h34234161_38234151,
        64'h3c234341_30234331,
        64'h34234321_38234291,
        64'h3c234481_3023bb01,
        64'h01138082_61657406,
        64'h70a6db7f_f0ef1828,
        64'h102cf29f_f0ef0028,
        64'h4681082c_1030e79f,
        64'hf0ef6027_b5030000,
        64'h0797e0be_4595603c,
        64'hfc3e4699_00b07c1c,
        64'h2f0000ef_f03e6c1c,
        64'hec3e681c_e83ef486,
        64'h00a8641c_e43e4661,
        64'h02040593_601c7064,
        64'h04130000_0417f0a2,
        64'h7159b7f9_f27ff0ef,
        64'h4511b7d1_f2fff0ef,
        64'h45058082_61054501,
        64'h64a26442_60e2eb7f,
        64'hf0ef45b1_46918622,
        64'hc3852781_4d3c66e7,
        64'hb5030000_07970007,
        64'h2023c78d_2781431c,
        64'h6807b703_00000797,
        64'hc3980007_a0234705,
        64'h6907b783_00000797,
        64'hf13ff0ef_45c18626,
        64'h46916a27_b5030000,
        64'h0797f25f_f0ef853e,
        64'h862a8432_45854691,
        64'h84ae10d7_a023e426,
        64'he822ec06_11016c67,
        64'hb7830000_07978082,
        64'h01410015_3513157d,
        64'h60a2fcbf_f0efe406,
        64'h1141b7fd_4501f06d,
        64'hfcbff0ef_347d8082,
        64'h01416402_60a2c789,
        64'h27815bbc_45057067,
        64'hb7830000_07976814,
        64'h0413e406_00989437,
        64'he0221141_bfdd2785,
        64'h00018082_00a7c363,
        64'h4781bfd1_060536fd,
        64'h2885c398_97aa97ae,
        64'h83f51782_411807bb,
        64'heb892701_0036f793,
        64'h8f5d0087_171b0006,
        64'h47838082_0006d363,
        64'hfff7881b_47014881,
        64'h36fd81f5_158202f6,
        64'hc7bb4791_b7d536fd,
        64'h06110107_a02397aa,
        64'h97ae83f5_00062803,
        64'h02069793_808200e6,
        64'h9363577d_36fd81f5,
        64'h1582b7ed_052136fd,
        64'hc38c97b2_83f90206,
        64'h9793410c_808200e6,
        64'h9363577d_952e36fd,
        64'h81f51582_8082c190,
        64'h95aa81f5_15828082,
        64'h418895aa_81f51582,
        64'hb7cd0006_0023b7e5,
        64'h00d60023_00d556b3,
        64'h0036969b_40e886bb,
        64'h00f6cb63_b7c50705,
        64'h01d60023_00d81663,
        64'h00e58633_bfc92000,
        64'h07938082_851a00de,
        64'h57630007_069bf800,
        64'h0e9388f2_87420077,
        64'h8e1b0107_87bbff83,
        64'h079b4037_581b4037,
        64'hd31b9f99_40000793,
        64'h02e7d963_1c000793,
        64'h1ff57713_80820015,
        64'h35138d1d_41dc4148,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00048067,
        64'h01f49493_0010049b,
        64'he3058593_00001597,
        64'hf1402573_ff2496e3,
        64'h00100493_0004a903,
        64'h04048493_01a49493,
        64'h0210049b_0924a4af,
        64'h00190913_04048493,
        64'h01a49493_0210049b,
        64'hff2496e3_f14024f3,
        64'h0004a903_04048493,
        64'h01a49493_0210049b,
        64'h055000ef_01a11113,
        64'h0210011b_01249863,
        64'hf1402973_00000493
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
